/home/pasam/common/Desktop/ECE581-2023/lab3-Chetanalahari-master/apr/work/saed32nm_hvt_1p9m.lef