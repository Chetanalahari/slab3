

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO ORCA_TOP 
  PIN sdram_clk 
    ANTENNAPARTIALMETALAREA 21.1396 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.377686 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0708 LAYER M6 ; 
    ANTENNAMAXAREACAR 309.929 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 5.58279 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.68306 LAYER VIA6 ;
  END sdram_clk
  PIN sys_2x_clk 
    ANTENNAPARTIALMETALAREA 9.38678 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.168038 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0579 LAYER M6 ; 
    ANTENNAMAXAREACAR 283.462 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 5.13132 LAYER M6 ;
    ANTENNAMAXCUTCAR 1.26582 LAYER VIA6 ;
  END sys_2x_clk
  PIN shutdown 
  END shutdown
  PIN test_mode 
    ANTENNAPARTIALMETALAREA 0.446648 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.016056 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1362 LAYER M6 ; 
    ANTENNAMAXAREACAR 59.436 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2.13143 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.556103 LAYER VIA6 ;
  END test_mode
  PIN test_si[5] 
    ANTENNAPARTIALMETALAREA 3.32421 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.118714 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 LAYER M6 ; 
    ANTENNAMAXAREACAR 211.306 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 7.55624 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.609573 LAYER VIA6 ;
  END test_si[5]
  PIN test_si[4] 
    ANTENNAPARTIALMETALAREA 2.12394 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.075944 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 LAYER M6 ; 
    ANTENNAMAXAREACAR 119.553 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 4.28667 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.609573 LAYER VIA6 ;
  END test_si[4]
  PIN test_si[3] 
    ANTENNAPARTIALMETALAREA 2.59218 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.09257 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1464 LAYER M6 ; 
    ANTENNAMAXAREACAR 18.9351 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 0.679003 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.0853825 LAYER VIA6 ;
  END test_si[3]
  PIN test_si[2] 
    ANTENNAPARTIALMETALAREA 0.43864 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.015658 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ; 
    ANTENNAMAXAREACAR 136.955 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 4.89276 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.595238 LAYER VIA6 ;
  END test_si[2]
  PIN test_si[1] 
    ANTENNAPARTIALMETALAREA 0.132208 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004714 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.051 LAYER M6 ; 
    ANTENNAMAXAREACAR 18.134 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 0.65851 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.348863 LAYER VIA6 ;
  END test_si[1]
  PIN test_si[0] 
    ANTENNAPARTIALMETALAREA 1.08555 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.038762 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ; 
    ANTENNAMAXAREACAR 95.6106 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 3.41619 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.595238 LAYER VIA6 ;
  END test_si[0]
  PIN test_so[5] 
    ANTENNADIFFAREA 0.6952 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.915312 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.032682 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0477 LAYER M6 ; 
    ANTENNAMAXAREACAR 109.794 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 3.92924 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.55313 LAYER VIA6 ;
  END test_so[5]
  PIN test_so[4] 
    ANTENNADIFFAREA 0.6952 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.064112 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.002282 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0477 LAYER M6 ; 
    ANTENNAMAXAREACAR 90.4723 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 3.24362 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.538467 LAYER VIA6 ;
  END test_so[4]
  PIN test_so[3] 
    ANTENNADIFFAREA 0.6952 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 7.93624 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.283526 LAYER M6 ;
  END test_so[3]
  PIN test_so[2] 
    ANTENNADIFFAREA 0.6952 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.302448 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.010794 LAYER M6 ;
  END test_so[2]
  PIN test_so[1] 
    ANTENNADIFFAREA 0.6952 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.132208 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004714 LAYER M6 ;
  END test_so[1]
  PIN test_so[0] 
    ANTENNADIFFAREA 0.6952 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.370544 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.013226 LAYER M6 ;
  END test_so[0]
  PIN scan_enable 
    ANTENNAPARTIALMETALAREA 0.302448 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.010794 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1464 LAYER M6 ; 
    ANTENNAMAXAREACAR 15.3303 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 0.55026 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.0853825 LAYER VIA6 ;
  END scan_enable
  PIN ate_clk 
    ANTENNAPARTIALMETALAREA 20.8362 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.372268 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0921 LAYER M6 ; 
    ANTENNAMAXAREACAR 252.304 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 4.54662 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.949367 LAYER VIA6 ;
  END ate_clk
  PIN occ_bypass 
  END occ_bypass
  PIN occ_reset 
  END occ_reset
  PIN pclk 
    ANTENNAPARTIALMETALAREA 7.34558 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.131364 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0579 LAYER M6 ; 
    ANTENNAMAXAREACAR 217.111 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 3.93995 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.949367 LAYER VIA6 ;
  END pclk
  PIN prst_n 
    ANTENNAPARTIALMETALAREA 0.140216 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.005112 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0471 LAYER M6 ; 
    ANTENNAMAXAREACAR 113.709 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 4.07326 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.550122 LAYER VIA6 ;
  END prst_n
  PIN pidsel 
  END pidsel
  PIN pgnt_n 
  END pgnt_n
  PIN pad_in[31] 
    ANTENNAPARTIALMETALAREA 1.25579 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.044842 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 LAYER M6 ; 
    ANTENNAMAXAREACAR 68.4903 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2.46316 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.534188 LAYER VIA6 ;
  END pad_in[31]
  PIN pad_in[30] 
    ANTENNAPARTIALMETALAREA 0.132208 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004714 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 LAYER M6 ; 
    ANTENNAMAXAREACAR 52.425 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1.8894 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.534188 LAYER VIA6 ;
  END pad_in[30]
  PIN pad_in[29] 
    ANTENNAPARTIALMETALAREA 1.08555 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.038762 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 LAYER M6 ; 
    ANTENNAMAXAREACAR 63.8212 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2.29641 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.534188 LAYER VIA6 ;
  END pad_in[29]
  PIN pad_in[28] 
    ANTENNAPARTIALMETALAREA 0.847216 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.03025 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 LAYER M6 ; 
    ANTENNAMAXAREACAR 59.8198 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2.1535 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.609573 LAYER VIA6 ;
  END pad_in[28]
  PIN pad_in[27] 
    ANTENNAPARTIALMETALAREA 0.030064 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.001066 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 LAYER M6 ; 
    ANTENNAMAXAREACAR 56.9569 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2.05128 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.534188 LAYER VIA6 ;
  END pad_in[27]
  PIN pad_in[26] 
    ANTENNAPARTIALMETALAREA 1.08555 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.038762 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 LAYER M6 ; 
    ANTENNAMAXAREACAR 52.4848 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1.89154 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.534188 LAYER VIA6 ;
  END pad_in[26]
  PIN pad_in[25] 
    ANTENNAPARTIALMETALAREA 1.25579 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.044842 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 LAYER M6 ; 
    ANTENNAMAXAREACAR 63.586 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2.28758 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.520833 LAYER VIA6 ;
  END pad_in[25]
  PIN pad_in[24] 
    ANTENNAPARTIALMETALAREA 1.28984 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.046058 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 LAYER M6 ; 
    ANTENNAMAXAREACAR 59.981 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2.15883 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.520833 LAYER VIA6 ;
  END pad_in[24]
  PIN pad_in[23] 
    ANTENNAPARTIALMETALAREA 0.540784 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.019306 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 LAYER M6 ; 
    ANTENNAMAXAREACAR 86.0578 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 3.0906 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.534188 LAYER VIA6 ;
  END pad_in[23]
  PIN pad_in[22] 
    ANTENNAPARTIALMETALAREA 0.030064 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.001066 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 LAYER M6 ; 
    ANTENNAMAXAREACAR 72.7956 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2.61692 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.534188 LAYER VIA6 ;
  END pad_in[22]
  PIN pad_in[21] 
    ANTENNAPARTIALMETALAREA 0.200304 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.007146 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 LAYER M6 ; 
    ANTENNAMAXAREACAR 69.1579 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2.48701 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.534188 LAYER VIA6 ;
  END pad_in[21]
  PIN pad_in[20] 
    ANTENNAPARTIALMETALAREA 0.200304 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.007146 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 LAYER M6 ; 
    ANTENNAMAXAREACAR 90.3128 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 3.24667 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.534188 LAYER VIA6 ;
  END pad_in[20]
  PIN pad_in[19] 
    ANTENNAPARTIALMETALAREA 0.813168 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.029034 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 LAYER M6 ; 
    ANTENNAMAXAREACAR 92.8622 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 3.33359 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.534188 LAYER VIA6 ;
  END pad_in[19]
  PIN pad_in[18] 
    ANTENNAPARTIALMETALAREA 0.09816 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.003498 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 LAYER M6 ; 
    ANTENNAMAXAREACAR 107.413 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 3.85325 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.534188 LAYER VIA6 ;
  END pad_in[18]
  PIN pad_in[17] 
    ANTENNAPARTIALMETALAREA 0.336496 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01201 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 LAYER M6 ; 
    ANTENNAMAXAREACAR 90.6797 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 3.25564 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.534188 LAYER VIA6 ;
  END pad_in[17]
  PIN pad_in[16] 
    ANTENNAPARTIALMETALAREA 0.302448 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.010794 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 LAYER M6 ; 
    ANTENNAMAXAREACAR 87.0421 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 3.12573 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.534188 LAYER VIA6 ;
  END pad_in[16]
  PIN pad_in[15] 
    ANTENNAPARTIALMETALAREA 0.030064 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.001066 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 LAYER M6 ; 
    ANTENNAMAXAREACAR 74.226 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2.66758 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.594333 LAYER VIA6 ;
  END pad_in[15]
  PIN pad_in[14] 
    ANTENNAPARTIALMETALAREA 0.09816 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.003498 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 LAYER M6 ; 
    ANTENNAMAXAREACAR 54.3647 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1.95825 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.594333 LAYER VIA6 ;
  END pad_in[14]
  PIN pad_in[13] 
    ANTENNAPARTIALMETALAREA 0.09816 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.003498 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 LAYER M6 ; 
    ANTENNAMAXAREACAR 65.4177 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2.353 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.594333 LAYER VIA6 ;
  END pad_in[13]
  PIN pad_in[12] 
    ANTENNAPARTIALMETALAREA 0.404592 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.014442 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 LAYER M6 ; 
    ANTENNAMAXAREACAR 65.301 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2.34883 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.594333 LAYER VIA6 ;
  END pad_in[12]
  PIN pad_in[11] 
    ANTENNAPARTIALMETALAREA 0.94936 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.033898 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 LAYER M6 ; 
    ANTENNAMAXAREACAR 87.7033 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 3.14892 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.520833 LAYER VIA6 ;
  END pad_in[11]
  PIN pad_in[10] 
    ANTENNAPARTIALMETALAREA 0.745072 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.026602 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 LAYER M6 ; 
    ANTENNAMAXAREACAR 80.9647 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2.90825 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.520833 LAYER VIA6 ;
  END pad_in[10]
  PIN pad_in[9] 
    ANTENNAPARTIALMETALAREA 0.60888 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.021738 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 LAYER M6 ; 
    ANTENNAMAXAREACAR 82.0287 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2.94625 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.520833 LAYER VIA6 ;
  END pad_in[9]
  PIN pad_in[8] 
    ANTENNAPARTIALMETALAREA 0.370544 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.013226 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 LAYER M6 ; 
    ANTENNAMAXAREACAR 74.7309 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2.69017 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.609573 LAYER VIA6 ;
  END pad_in[8]
  PIN pad_in[7] 
    ANTENNAPARTIALMETALAREA 0.302448 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.010794 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 LAYER M6 ; 
    ANTENNAMAXAREACAR 47.9807 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1.73025 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.594333 LAYER VIA6 ;
  END pad_in[7]
  PIN pad_in[6] 
    ANTENNAPARTIALMETALAREA 1.08555 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.038762 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 LAYER M6 ; 
    ANTENNAMAXAREACAR 51.6317 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1.86067 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.594333 LAYER VIA6 ;
  END pad_in[6]
  PIN pad_in[5] 
    ANTENNAPARTIALMETALAREA 0.43864 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.015658 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 LAYER M6 ; 
    ANTENNAMAXAREACAR 60.9113 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2.19208 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.594333 LAYER VIA6 ;
  END pad_in[5]
  PIN pad_in[4] 
    ANTENNAPARTIALMETALAREA 0.234352 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.008362 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 LAYER M6 ; 
    ANTENNAMAXAREACAR 48.2267 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1.73949 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.609573 LAYER VIA6 ;
  END pad_in[4]
  PIN pad_in[3] 
    ANTENNAPARTIALMETALAREA 0.745072 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.026602 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 LAYER M6 ; 
    ANTENNAMAXAREACAR 47.452 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1.71179 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.609573 LAYER VIA6 ;
  END pad_in[3]
  PIN pad_in[2] 
    ANTENNAPARTIALMETALAREA 0.540784 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.019306 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 LAYER M6 ; 
    ANTENNAMAXAREACAR 51.7573 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1.86556 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.609573 LAYER VIA6 ;
  END pad_in[2]
  PIN pad_in[1] 
    ANTENNAPARTIALMETALAREA 0.506736 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01809 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 LAYER M6 ; 
    ANTENNAMAXAREACAR 42.6632 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1.54077 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.609573 LAYER VIA6 ;
  END pad_in[1]
  PIN pad_in[0] 
    ANTENNAPARTIALMETALAREA 0.813168 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.029034 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 LAYER M6 ; 
    ANTENNAMAXAREACAR 42.6607 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1.54025 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.520833 LAYER VIA6 ;
  END pad_in[0]
  PIN pad_out[31] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.200304 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.007146 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ; 
    ANTENNAMAXAREACAR 116.36 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 4.17067 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.714286 LAYER VIA6 ;
  END pad_out[31]
  PIN pad_out[30] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.132208 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004714 LAYER M6 ;
  END pad_out[30]
  PIN pad_out[29] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.09816 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.003498 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ; 
    ANTENNAMAXAREACAR 134.398 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 4.81029 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.714286 LAYER VIA6 ;
  END pad_out[29]
  PIN pad_out[28] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.132208 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004714 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ; 
    ANTENNAMAXAREACAR 33.3717 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1.198 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.595238 LAYER VIA6 ;
  END pad_out[28]
  PIN pad_out[27] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.302448 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.010794 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ; 
    ANTENNAMAXAREACAR 174.308 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 6.23143 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.595238 LAYER VIA6 ;
  END pad_out[27]
  PIN pad_out[26] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.030064 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.001066 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ; 
    ANTENNAMAXAREACAR 94.235 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 3.37629 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.595238 LAYER VIA6 ;
  END pad_out[26]
  PIN pad_out[25] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.064112 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.002282 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ; 
    ANTENNAMAXAREACAR 76.9652 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 2.75914 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.595238 LAYER VIA6 ;
  END pad_out[25]
  PIN pad_out[24] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.09816 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.003498 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ; 
    ANTENNAMAXAREACAR 94.9264 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 3.40095 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.595238 LAYER VIA6 ;
  END pad_out[24]
  PIN pad_out[23] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.2684 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.009578 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ; 
    ANTENNAMAXAREACAR 218.172 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 7.79762 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.595238 LAYER VIA6 ;
  END pad_out[23]
  PIN pad_out[22] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.030064 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.001066 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ; 
    ANTENNAMAXAREACAR 87.1618 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 3.11905 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.595238 LAYER VIA6 ;
  END pad_out[22]
  PIN pad_out[21] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.030064 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.001066 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ; 
    ANTENNAMAXAREACAR 154.873 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 5.53695 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.595238 LAYER VIA6 ;
  END pad_out[21]
  PIN pad_out[20] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.404592 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.014442 LAYER M6 ;
  END pad_out[20]
  PIN pad_out[19] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.132208 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004714 LAYER M6 ;
  END pad_out[19]
  PIN pad_out[18] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.200304 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.007146 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ; 
    ANTENNAMAXAREACAR 116.433 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 4.1641 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.595238 LAYER VIA6 ;
  END pad_out[18]
  PIN pad_out[17] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 1.53809 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.054924 LAYER M6 ;
  END pad_out[17]
  PIN pad_out[16] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.506736 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01809 LAYER M6 ;
  END pad_out[16]
  PIN pad_out[15] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.064112 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.002282 LAYER M6 ;
  END pad_out[15]
  PIN pad_out[14] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.2684 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.009578 LAYER M6 ;
  END pad_out[14]
  PIN pad_out[13] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 1.36785 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.048844 LAYER M6 ;
  END pad_out[13]
  PIN pad_out[12] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.09816 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.003498 LAYER M6 ;
  END pad_out[12]
  PIN pad_out[11] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 1.53809 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.054924 LAYER M6 ;
  END pad_out[11]
  PIN pad_out[10] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 1.08555 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.038762 LAYER M6 ;
  END pad_out[10]
  PIN pad_out[9] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.030064 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.001066 LAYER M6 ;
  END pad_out[9]
  PIN pad_out[8] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.200304 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.007146 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 LAYER M6 ; 
    ANTENNAMAXAREACAR 54.1473 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 1.94419 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.595238 LAYER VIA6 ;
  END pad_out[8]
  PIN pad_out[7] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.234352 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.008362 LAYER M6 ;
  END pad_out[7]
  PIN pad_out[6] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.064112 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.002282 LAYER M6 ;
  END pad_out[6]
  PIN pad_out[5] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 1.94526 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.069466 LAYER M6 ;
  END pad_out[5]
  PIN pad_out[4] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.2684 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.009578 LAYER M6 ;
  END pad_out[4]
  PIN pad_out[3] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 1.08555 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.038762 LAYER M6 ;
  END pad_out[3]
  PIN pad_out[2] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 1.0515 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.037546 LAYER M6 ;
  END pad_out[2]
  PIN pad_out[1] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 1.59627 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.057002 LAYER M6 ;
  END pad_out[1]
  PIN pad_out[0] 
    ANTENNADIFFAREA 2.4808 LAYER M6 ; 
    ANTENNAPARTIALMETALAREA 0.030064 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.001066 LAYER M6 ;
  END pad_out[0]
  PIN ppar_in 
  END ppar_in
  PIN pc_be_in[3] 
    ANTENNAPARTIALMETALAREA 0.676976 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.02417 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1401 LAYER M6 ; 
    ANTENNAMAXAREACAR 14.0775 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 0.507829 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.322652 LAYER VIA6 ;
  END pc_be_in[3]
  PIN pc_be_in[2] 
    ANTENNAPARTIALMETALAREA 0.60888 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.021738 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1122 LAYER M6 ; 
    ANTENNAMAXAREACAR 10.9005 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 0.389854 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.290734 LAYER VIA6 ;
  END pc_be_in[2]
  PIN pc_be_in[1] 
    ANTENNAPARTIALMETALAREA 0.574832 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.020522 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1122 LAYER M6 ; 
    ANTENNAMAXAREACAR 10.1828 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 0.363747 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.271349 LAYER VIA6 ;
  END pc_be_in[1]
  PIN pc_be_in[0] 
    ANTENNAPARTIALMETALAREA 0.676976 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.02417 LAYER M6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1401 LAYER M6 ; 
    ANTENNAMAXAREACAR 13.0744 LAYER M6 ;
    ANTENNAMAXSIDEAREACAR 0.470839 LAYER M6 ;
    ANTENNAMAXCUTCAR 0.265328 LAYER VIA6 ;
  END pc_be_in[0]
  PIN pframe_n_in 
  END pframe_n_in
  PIN ptrdy_n_in 
  END ptrdy_n_in
  PIN pirdy_n_in 
  END pirdy_n_in
  PIN pdevsel_n_in 
  END pdevsel_n_in
  PIN pstop_n_in 
  END pstop_n_in
  PIN pperr_n_in 
  END pperr_n_in
  PIN pserr_n_in 
  END pserr_n_in
  PIN pm66en 
  END pm66en
  PIN sd_A[9] 
    ANTENNADIFFAREA 0.3976 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.200304 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.007146 LAYER M8 ;
  END sd_A[9]
  PIN sd_A[8] 
    ANTENNADIFFAREA 0.3976 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.472688 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.016874 LAYER M8 ;
  END sd_A[8]
  PIN sd_A[7] 
    ANTENNADIFFAREA 0.2488 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.404592 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.014442 LAYER M8 ;
  END sd_A[7]
  PIN sd_A[6] 
    ANTENNADIFFAREA 0.2488 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.00044 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 8e-06 LAYER M8 ;
  END sd_A[6]
  PIN sd_A[5] 
    ANTENNAPARTIALMETALAREA 0.154608 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.005024 LAYER M8 ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA8 ;
    ANTENNADIFFAREA 0.3976 LAYER M9 ; 
    ANTENNAPARTIALMETALAREA 0.22496 LAYER M9 ;
    ANTENNAPARTIALMETALSIDEAREA 0.003132 LAYER M9 ;
  END sd_A[5]
  PIN sd_A[4] 
    ANTENNAPARTIALMETALAREA 0.094512 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.002982 LAYER M8 ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA8 ;
    ANTENNADIFFAREA 0.3976 LAYER M9 ; 
    ANTENNAPARTIALMETALAREA 2.68128 LAYER M9 ;
    ANTENNAPARTIALMETALSIDEAREA 0.033836 LAYER M9 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 LAYER M9 ; 
    ANTENNAMAXAREACAR 181.726 LAYER M9 ;
    ANTENNAMAXSIDEAREACAR 3.53343 LAYER M9 ;
    ANTENNAMAXCUTCAR 1.6381 LAYER VIARDL ;
  END sd_A[4]
  PIN sd_A[3] 
    ANTENNADIFFAREA 0.3976 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.540784 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.019306 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ; 
    ANTENNAMAXAREACAR 97.8532 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 3.50971 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.833333 LAYER VIA8 ;
  END sd_A[3]
  PIN sd_A[2] 
    ANTENNADIFFAREA 0.3976 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.2684 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.009578 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 LAYER M8 ; 
    ANTENNAMAXAREACAR 143.651 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 5.14533 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.833333 LAYER VIA8 ;
  END sd_A[2]
  PIN sd_A[1] 
    ANTENNADIFFAREA 0.3976 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.200304 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.007146 LAYER M8 ;
  END sd_A[1]
  PIN sd_A[0] 
    ANTENNAPARTIALMETALAREA 0.563184 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.019616 LAYER M8 ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA8 ;
    ANTENNADIFFAREA 0.3976 LAYER M9 ; 
    ANTENNAPARTIALMETALAREA 0.54112 LAYER M9 ;
    ANTENNAPARTIALMETALSIDEAREA 0.007084 LAYER M9 ;
  END sd_A[0]
  PIN sd_CK 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.132208 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004714 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.822 LAYER M8 ; 
    ANTENNAMAXAREACAR 144.524 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 5.17062 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.51949 LAYER VIA8 ;
  END sd_CK
  PIN sd_CKn 
    ANTENNADIFFAREA 1.2904 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.064112 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.002282 LAYER M8 ;
  END sd_CKn
  PIN sd_LD 
    ANTENNADIFFAREA 0.2488 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.472688 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.016874 LAYER M8 ;
  END sd_LD
  PIN sd_RW 
    ANTENNAPARTIALMETALAREA 0.774512 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.02726 LAYER M8 ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA8 ;
    ANTENNADIFFAREA 0.2488 LAYER M9 ; 
    ANTENNAPARTIALMETALAREA 0.24928 LAYER M9 ;
    ANTENNAPARTIALMETALSIDEAREA 0.003436 LAYER M9 ;
  END sd_RW
  PIN sd_BWS[1] 
    ANTENNADIFFAREA 0.3976 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.132208 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004714 LAYER M8 ;
  END sd_BWS[1]
  PIN sd_BWS[0] 
    ANTENNADIFFAREA 0.2488 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.684016 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.024518 LAYER M8 ;
  END sd_BWS[0]
  PIN sd_DQ_in[31] 
    ANTENNAPARTIALMETALAREA 0.9788 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.034556 LAYER M8 ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA8 ;
    ANTENNAPARTIALMETALAREA 0.5168 LAYER M9 ;
    ANTENNAPARTIALMETALSIDEAREA 0.00678 LAYER M9 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M9 ; 
    ANTENNAMAXAREACAR 90.6249 LAYER M9 ;
    ANTENNAMAXSIDEAREACAR 2.74979 LAYER M9 ;
    ANTENNAMAXCUTCAR 1.52591 LAYER VIARDL ;
  END sd_DQ_in[31]
  PIN sd_DQ_in[30] 
    ANTENNAPARTIALMETALAREA 0.480696 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.017272 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 39.4198 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 1.43477 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.738397 LAYER VIA8 ;
  END sd_DQ_in[30]
  PIN sd_DQ_in[29] 
    ANTENNAPARTIALMETALAREA 1.46809 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.052536 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 121.261 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 4.35764 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.812827 LAYER VIA8 ;
  END sd_DQ_in[29]
  PIN sd_DQ_in[28] 
    ANTENNAPARTIALMETALAREA 0.336496 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01201 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 36.5213 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 1.3265 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.812827 LAYER VIA8 ;
  END sd_DQ_in[28]
  PIN sd_DQ_in[27] 
    ANTENNAPARTIALMETALAREA 0.07212 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.00268 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 125.423 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 4.50633 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.738397 LAYER VIA8 ;
  END sd_DQ_in[27]
  PIN sd_DQ_in[26] 
    ANTENNAPARTIALMETALAREA 1.10207 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.039464 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 162.923 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 5.84557 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.812827 LAYER VIA8 ;
  END sd_DQ_in[26]
  PIN sd_DQ_in[25] 
    ANTENNAPARTIALMETALAREA 1.39198 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.049706 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 66.9017 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 2.41156 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.812827 LAYER VIA8 ;
  END sd_DQ_in[25]
  PIN sd_DQ_in[24] 
    ANTENNAPARTIALMETALAREA 1.25572 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.044936 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 209.737 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 7.51688 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.738397 LAYER VIA8 ;
  END sd_DQ_in[24]
  PIN sd_DQ_in[23] 
    ANTENNAPARTIALMETALAREA 0.540784 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.019306 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 45.5002 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 1.64717 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.738397 LAYER VIA8 ;
  END sd_DQ_in[23]
  PIN sd_DQ_in[22] 
    ANTENNAPARTIALMETALAREA 0.315496 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01077 LAYER M8 ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA8 ;
    ANTENNAPARTIALMETALAREA 0.80864 LAYER M9 ;
    ANTENNAPARTIALMETALSIDEAREA 0.010428 LAYER M9 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M9 ; 
    ANTENNAMAXAREACAR 109.404 LAYER M9 ;
    ANTENNAMAXSIDEAREACAR 3.1346 LAYER M9 ;
    ANTENNAMAXCUTCAR 1.52591 LAYER VIARDL ;
  END sd_DQ_in[22]
  PIN sd_DQ_in[21] 
    ANTENNAPARTIALMETALAREA 0.132208 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004714 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 43.3452 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 1.57021 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.738397 LAYER VIA8 ;
  END sd_DQ_in[21]
  PIN sd_DQ_in[20] 
    ANTENNAPARTIALMETALAREA 0.218728 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.007804 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 186.649 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 6.68819 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.738397 LAYER VIA8 ;
  END sd_DQ_in[20]
  PIN sd_DQ_in[19] 
    ANTENNAPARTIALMETALAREA 0.00044 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 8e-06 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 44.6306 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 1.61612 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.738397 LAYER VIA8 ;
  END sd_DQ_in[19]
  PIN sd_DQ_in[18] 
    ANTENNAPARTIALMETALAREA 0.140216 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.005112 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 109.676 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 3.94802 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.738397 LAYER VIA8 ;
  END sd_DQ_in[18]
  PIN sd_DQ_in[17] 
    ANTENNAPARTIALMETALAREA 0.981432 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.035252 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 123.713 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 4.44928 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.812827 LAYER VIA8 ;
  END sd_DQ_in[17]
  PIN sd_DQ_in[16] 
    ANTENNAPARTIALMETALAREA 0.426992 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.014752 LAYER M8 ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA8 ;
    ANTENNAPARTIALMETALAREA 9 LAYER M9 ;
    ANTENNAPARTIALMETALSIDEAREA 0.012 LAYER M9 ;
    ANTENNAPARTIALCUTAREA 4 LAYER VIARDL ;
    ANTENNAPARTIALMETALAREA 31.456 LAYER MRDL ;
    ANTENNAPARTIALMETALSIDEAREA 0.033456 LAYER MRDL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER MRDL ; 
    ANTENNAMAXAREACAR 1734.88 LAYER MRDL ;
    ANTENNAMAXSIDEAREACAR 2.91941 LAYER MRDL ;
  END sd_DQ_in[16]
  PIN sd_DQ_in[15] 
    ANTENNAPARTIALMETALAREA 0.200304 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.007146 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 174.434 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 6.25603 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.738397 LAYER VIA8 ;
  END sd_DQ_in[15]
  PIN sd_DQ_in[14] 
    ANTENNAPARTIALMETALAREA 1.10795 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.039072 LAYER M8 ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA8 ;
    ANTENNAPARTIALMETALAREA 0.152 LAYER M9 ;
    ANTENNAPARTIALMETALSIDEAREA 0.00222 LAYER M9 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M9 ; 
    ANTENNAMAXAREACAR 75.8887 LAYER M9 ;
    ANTENNAMAXSIDEAREACAR 2.58489 LAYER M9 ;
    ANTENNAMAXCUTCAR 1.52591 LAYER VIARDL ;
  END sd_DQ_in[14]
  PIN sd_DQ_in[13] 
    ANTENNAPARTIALMETALAREA 1.66437 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.059434 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0732 LAYER M8 ; 
    ANTENNAMAXAREACAR 45.7183 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 1.64005 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.287268 LAYER VIA8 ;
  END sd_DQ_in[13]
  PIN sd_DQ_in[12] 
    ANTENNAPARTIALMETALAREA 0.889272 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.031864 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 250.557 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 8.97536 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.812827 LAYER VIA8 ;
  END sd_DQ_in[12]
  PIN sd_DQ_in[11] 
    ANTENNAPARTIALMETALAREA 0.07212 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.00268 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 34.1381 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 1.24616 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.738397 LAYER VIA8 ;
  END sd_DQ_in[11]
  PIN sd_DQ_in[10] 
    ANTENNAPARTIALMETALAREA 0.85112 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.029996 LAYER M8 ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA8 ;
    ANTENNAPARTIALMETALAREA 0.61408 LAYER M9 ;
    ANTENNAPARTIALMETALSIDEAREA 0.007996 LAYER M9 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M9 ; 
    ANTENNAMAXAREACAR 93.2929 LAYER M9 ;
    ANTENNAMAXSIDEAREACAR 2.74979 LAYER M9 ;
    ANTENNAMAXCUTCAR 1.52591 LAYER VIARDL ;
  END sd_DQ_in[10]
  PIN sd_DQ_in[9] 
    ANTENNAPARTIALMETALAREA 1.46809 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.052536 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 87.141 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 3.13907 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.738397 LAYER VIA8 ;
  END sd_DQ_in[9]
  PIN sd_DQ_in[8] 
    ANTENNAPARTIALMETALAREA 0.676976 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.02417 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 40.5186 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 1.46928 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.812827 LAYER VIA8 ;
  END sd_DQ_in[8]
  PIN sd_DQ_in[7] 
    ANTENNAPARTIALMETALAREA 0.813168 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.029034 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 250.219 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 8.95857 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.738397 LAYER VIA8 ;
  END sd_DQ_in[7]
  PIN sd_DQ_in[6] 
    ANTENNAPARTIALMETALAREA 0.472688 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.016874 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 60.6998 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 2.19409 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.738397 LAYER VIA8 ;
  END sd_DQ_in[6]
  PIN sd_DQ_in[5] 
    ANTENNAPARTIALMETALAREA 1.56222 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.055786 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2928 LAYER M8 ; 
    ANTENNAMAXAREACAR 8.93131 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 0.321455 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.0597678 LAYER VIA8 ;
  END sd_DQ_in[5]
  PIN sd_DQ_in[4] 
    ANTENNAPARTIALMETALAREA 0.557304 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.020008 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 200.275 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 7.17958 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.812827 LAYER VIA8 ;
  END sd_DQ_in[4]
  PIN sd_DQ_in[3] 
    ANTENNAPARTIALMETALAREA 0.00044 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 8e-06 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 163.293 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 5.85814 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.738397 LAYER VIA8 ;
  END sd_DQ_in[3]
  PIN sd_DQ_in[2] 
    ANTENNAPARTIALMETALAREA 0.2684 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.009578 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 159.409 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 5.71941 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.738397 LAYER VIA8 ;
  END sd_DQ_in[2]
  PIN sd_DQ_in[1] 
    ANTENNAPARTIALMETALAREA 0.763496 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.02726 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 54.6438 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 1.97376 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.738397 LAYER VIA8 ;
  END sd_DQ_in[1]
  PIN sd_DQ_in[0] 
    ANTENNAPARTIALMETALAREA 0.94936 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.033898 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 53.5663 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 1.93527 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.812827 LAYER VIA8 ;
  END sd_DQ_in[0]
  PIN sd_DQ_out[31] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.064112 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.002282 LAYER M8 ;
  END sd_DQ_out[31]
  PIN sd_DQ_out[30] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.404592 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.014442 LAYER M8 ;
  END sd_DQ_out[30]
  PIN sd_DQ_out[29] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.064112 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.002282 LAYER M8 ;
  END sd_DQ_out[29]
  PIN sd_DQ_out[28] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.132208 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004714 LAYER M8 ;
  END sd_DQ_out[28]
  PIN sd_DQ_out[27] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.404592 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.014442 LAYER M8 ;
  END sd_DQ_out[27]
  PIN sd_DQ_out[26] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.064112 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.002282 LAYER M8 ;
  END sd_DQ_out[26]
  PIN sd_DQ_out[25] 
    ANTENNADIFFAREA 0.3976 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.200304 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.007146 LAYER M8 ;
  END sd_DQ_out[25]
  PIN sd_DQ_out[24] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.132208 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004714 LAYER M8 ;
  END sd_DQ_out[24]
  PIN sd_DQ_out[23] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.336496 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01201 LAYER M8 ;
  END sd_DQ_out[23]
  PIN sd_DQ_out[22] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.132208 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004714 LAYER M8 ;
  END sd_DQ_out[22]
  PIN sd_DQ_out[21] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.2684 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.009578 LAYER M8 ;
  END sd_DQ_out[21]
  PIN sd_DQ_out[20] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.336496 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01201 LAYER M8 ;
  END sd_DQ_out[20]
  PIN sd_DQ_out[19] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.404592 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.014442 LAYER M8 ;
  END sd_DQ_out[19]
  PIN sd_DQ_out[18] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.2684 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.009578 LAYER M8 ;
  END sd_DQ_out[18]
  PIN sd_DQ_out[17] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.064112 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.002282 LAYER M8 ;
  END sd_DQ_out[17]
  PIN sd_DQ_out[16] 
    ANTENNADIFFAREA 0.3976 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.200304 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.007146 LAYER M8 ;
  END sd_DQ_out[16]
  PIN sd_DQ_out[15] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.132208 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004714 LAYER M8 ;
  END sd_DQ_out[15]
  PIN sd_DQ_out[14] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.064112 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.002282 LAYER M8 ;
  END sd_DQ_out[14]
  PIN sd_DQ_out[13] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.2684 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.009578 LAYER M8 ;
  END sd_DQ_out[13]
  PIN sd_DQ_out[12] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.336496 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01201 LAYER M8 ;
  END sd_DQ_out[12]
  PIN sd_DQ_out[11] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.064112 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.002282 LAYER M8 ;
  END sd_DQ_out[11]
  PIN sd_DQ_out[10] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.2684 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.009578 LAYER M8 ;
  END sd_DQ_out[10]
  PIN sd_DQ_out[9] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.132208 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004714 LAYER M8 ;
  END sd_DQ_out[9]
  PIN sd_DQ_out[8] 
    ANTENNADIFFAREA 0.3976 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.200304 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.007146 LAYER M8 ;
  END sd_DQ_out[8]
  PIN sd_DQ_out[7] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.064112 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.002282 LAYER M8 ;
  END sd_DQ_out[7]
  PIN sd_DQ_out[6] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.132208 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004714 LAYER M8 ;
  END sd_DQ_out[6]
  PIN sd_DQ_out[5] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.064112 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.002282 LAYER M8 ;
  END sd_DQ_out[5]
  PIN sd_DQ_out[4] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.200304 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.007146 LAYER M8 ;
  END sd_DQ_out[4]
  PIN sd_DQ_out[3] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.00044 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 8e-06 LAYER M8 ;
  END sd_DQ_out[3]
  PIN sd_DQ_out[2] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.2684 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.009578 LAYER M8 ;
  END sd_DQ_out[2]
  PIN sd_DQ_out[1] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.404592 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.014442 LAYER M8 ;
  END sd_DQ_out[1]
  PIN sd_DQ_out[0] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.064112 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.002282 LAYER M8 ;
  END sd_DQ_out[0]
  PIN sd_DQ_en[29] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.311184 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.011106 LAYER M8 ;
  END sd_DQ_en[29]
  PIN sd_DQ_en[30] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.31432 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01133 LAYER M8 ;
  END sd_DQ_en[30]
  PIN sd_DQ_en[31] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.312752 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.011274 LAYER M8 ;
  END sd_DQ_en[31]
  PIN sd_DQ_en[23] 
    ANTENNADIFFAREA 1.2904 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.988224 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.035286 LAYER M8 ;
  END sd_DQ_en[23]
  PIN sd_DQ_en[24] 
    ANTENNADIFFAREA 1.2904 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.99136 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.03551 LAYER M8 ;
  END sd_DQ_en[24]
  PIN sd_DQ_en[25] 
    ANTENNADIFFAREA 1.2904 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.99136 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.03551 LAYER M8 ;
  END sd_DQ_en[25]
  PIN sd_DQ_en[26] 
    ANTENNADIFFAREA 1.2904 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.99136 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.03551 LAYER M8 ;
  END sd_DQ_en[26]
  PIN sd_DQ_en[27] 
    ANTENNADIFFAREA 1.2904 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.99136 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.03551 LAYER M8 ;
  END sd_DQ_en[27]
  PIN sd_DQ_en[28] 
    ANTENNADIFFAREA 1.2904 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.989792 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.035454 LAYER M8 ;
  END sd_DQ_en[28]
  PIN sd_DQ_en[16] 
    ANTENNADIFFAREA 1.2904 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.47144 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.017038 LAYER M8 ;
  END sd_DQ_en[16]
  PIN sd_DQ_en[18] 
    ANTENNADIFFAREA 1.2904 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.479448 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.017436 LAYER M8 ;
  END sd_DQ_en[18]
  PIN sd_DQ_en[20] 
    ANTENNADIFFAREA 1.2904 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.480232 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.017492 LAYER M8 ;
  END sd_DQ_en[20]
  PIN sd_DQ_en[21] 
    ANTENNADIFFAREA 1.2904 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.474576 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.017262 LAYER M8 ;
  END sd_DQ_en[21]
  PIN sd_DQ_en[22] 
    ANTENNADIFFAREA 1.2904 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.473008 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.017206 LAYER M8 ;
  END sd_DQ_en[22]
  PIN sd_DQ_en[14] 
    ANTENNADIFFAREA 0.3976 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.472688 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.016874 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1098 LAYER M8 ; 
    ANTENNAMAXAREACAR 7.153 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 0.260528 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.159381 LAYER VIA8 ;
  END sd_DQ_en[14]
  PIN sd_DQ_en[12] 
    ANTENNADIFFAREA 0.3976 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.1536 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.005478 LAYER M8 ;
  END sd_DQ_en[12]
  PIN sd_DQ_en[13] 
    ANTENNADIFFAREA 0.3976 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.155168 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.005646 LAYER M8 ;
  END sd_DQ_en[13]
  PIN sd_DQ_en[10] 
    ANTENNADIFFAREA 1.2904 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.289008 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.010426 LAYER M8 ;
  END sd_DQ_en[10]
  PIN sd_DQ_en[11] 
    ANTENNADIFFAREA 1.2904 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.28744 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01037 LAYER M8 ;
  END sd_DQ_en[11]
  PIN sd_DQ_en[7] 
    ANTENNADIFFAREA 1.2904 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.285872 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.010202 LAYER M8 ;
  END sd_DQ_en[7]
  PIN sd_DQ_en[8] 
    ANTENNADIFFAREA 1.2904 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.289008 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.010426 LAYER M8 ;
  END sd_DQ_en[8]
  PIN sd_DQ_en[9] 
    ANTENNADIFFAREA 1.2904 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.289008 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.010426 LAYER M8 ;
  END sd_DQ_en[9]
  PIN sd_DQ_en[6] 
    ANTENNADIFFAREA 0.3976 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.132208 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004714 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1098 LAYER M8 ; 
    ANTENNAMAXAREACAR 9.62301 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 0.349617 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.182149 LAYER VIA8 ;
  END sd_DQ_en[6]
  PIN sd_DQ_en[1] 
    ANTENNADIFFAREA 1.2904 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.422064 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.015066 LAYER M8 ;
  END sd_DQ_en[1]
  PIN sd_DQ_en[2] 
    ANTENNADIFFAREA 1.2904 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.4252 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01529 LAYER M8 ;
  END sd_DQ_en[2]
  PIN sd_DQ_en[3] 
    ANTENNADIFFAREA 1.2904 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.4252 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01529 LAYER M8 ;
  END sd_DQ_en[3]
  PIN sd_DQ_en[4] 
    ANTENNADIFFAREA 1.2904 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.4252 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01529 LAYER M8 ;
  END sd_DQ_en[4]
  PIN sd_DQ_en[5] 
    ANTENNADIFFAREA 1.2904 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.423632 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.015234 LAYER M8 ;
  END sd_DQ_en[5]
  PIN sd_DQ_en[0] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.240824 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.008906 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ; 
    ANTENNAMAXAREACAR 6.57989 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 0.243333 LAYER M8 ;
  END sd_DQ_en[0]
  PIN sd_DQ_en[15] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.248832 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.009304 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ; 
    ANTENNAMAXAREACAR 6.79869 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 0.254208 LAYER M8 ;
  END sd_DQ_en[15]
  PIN sd_DQ_en[17] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.248832 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.009304 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ; 
    ANTENNAMAXAREACAR 38.5315 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 1.40022 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.68306 LAYER VIA8 ;
  END sd_DQ_en[17]
  PIN sd_DQ_en[19] 
    ANTENNADIFFAREA 0.6952 LAYER M8 ; 
    ANTENNAPARTIALMETALAREA 0.246984 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.009238 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 LAYER M8 ; 
    ANTENNAMAXAREACAR 6.7482 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 0.252404 LAYER M8 ;
  END sd_DQ_en[19]
  PIN pll_bypass 
    ANTENNAPARTIALMETALAREA 0.480696 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.017272 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2478 LAYER M8 ; 
    ANTENNAMAXAREACAR 45.3915 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 1.63751 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.642212 LAYER VIA8 ;
  END pll_bypass
  PIN pll_reset 
    ANTENNAPARTIALMETALAREA 0.0066 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.00034 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 LAYER M8 ; 
    ANTENNAMAXAREACAR 42.7822 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 1.55485 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.812827 LAYER VIA8 ;
  END pll_reset
  PIN test_si7 
    ANTENNAPARTIALMETALAREA 0.276912 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.009882 LAYER M8 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0285 LAYER M8 ; 
    ANTENNAMAXAREACAR 435.416 LAYER M8 ;
    ANTENNAMAXSIDEAREACAR 15.5585 LAYER M8 ;
    ANTENNAMAXCUTCAR 0.67593 LAYER VIA8 ;
  END test_si7
  PIN test_so7 
    ANTENNAPARTIALMETALAREA 0.154608 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 0.005024 LAYER M8 ;
    ANTENNAPARTIALCUTAREA 0.0169 LAYER VIA8 ;
    ANTENNADIFFAREA 0.3976 LAYER M9 ; 
    ANTENNAPARTIALMETALAREA 0.37088 LAYER M9 ;
    ANTENNAPARTIALMETALSIDEAREA 0.004956 LAYER M9 ;
  END test_so7
END ORCA_TOP

END LIBRARY
