/home/pasam/common/Desktop/ECE581-2023/lab3-Chetanalahari-master/cadence_cap_tech/tech.lef